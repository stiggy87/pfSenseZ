`timescale 1 ps / 1 ps
// lib IP_Integrator_Lib
module pfSenseZ_wrapper
   (DDR_addr,
    DDR_ba,
    DDR_cas_n,
    DDR_ck_n,
    DDR_ck_p,
    DDR_cke,
    DDR_cs_n,
    DDR_dm,
    DDR_dq,
    DDR_dqs_n,
    DDR_dqs_p,
    DDR_odt,
    DDR_ras_n,
    DDR_reset_n,
    DDR_we_n,
    FIXED_IO_ddr_vrn,
    FIXED_IO_ddr_vrp,
    FIXED_IO_mio,
    FIXED_IO_ps_clk,
    FIXED_IO_ps_porb,
    FIXED_IO_ps_srstb,
    GMII_ETHERNET_1_col,
    GMII_ETHERNET_1_crs,
    GMII_ETHERNET_1_rx_clk,
    GMII_ETHERNET_1_rx_dv,
    GMII_ETHERNET_1_rx_er,
    GMII_ETHERNET_1_rxd,
    GMII_ETHERNET_1_tx_clk,
    GMII_ETHERNET_1_tx_en,
    GMII_ETHERNET_1_tx_er,
    GMII_ETHERNET_1_txd,
    btns_5bits_tri_io,
    leds_8bits_tri_o);
  inout [14:0]DDR_addr;
  inout [2:0]DDR_ba;
  inout DDR_cas_n;
  inout DDR_ck_n;
  inout DDR_ck_p;
  inout DDR_cke;
  inout DDR_cs_n;
  inout [3:0]DDR_dm;
  inout [31:0]DDR_dq;
  inout [3:0]DDR_dqs_n;
  inout [3:0]DDR_dqs_p;
  inout DDR_odt;
  inout DDR_ras_n;
  inout DDR_reset_n;
  inout DDR_we_n;
  inout FIXED_IO_ddr_vrn;
  inout FIXED_IO_ddr_vrp;
  inout [53:0]FIXED_IO_mio;
  inout FIXED_IO_ps_clk;
  inout FIXED_IO_ps_porb;
  inout FIXED_IO_ps_srstb;
  input GMII_ETHERNET_1_col;
  input GMII_ETHERNET_1_crs;
  input GMII_ETHERNET_1_rx_clk;
  input GMII_ETHERNET_1_rx_dv;
  input GMII_ETHERNET_1_rx_er;
  input [7:0]GMII_ETHERNET_1_rxd;
  input GMII_ETHERNET_1_tx_clk;
  output [0:0]GMII_ETHERNET_1_tx_en;
  output [0:0]GMII_ETHERNET_1_tx_er;
  output [7:0]GMII_ETHERNET_1_txd;
  inout [4:0]btns_5bits_tri_io;
  output [7:0]leds_8bits_tri_o;

  wire [14:0]DDR_addr;
  wire [2:0]DDR_ba;
  wire DDR_cas_n;
  wire DDR_ck_n;
  wire DDR_ck_p;
  wire DDR_cke;
  wire DDR_cs_n;
  wire [3:0]DDR_dm;
  wire [31:0]DDR_dq;
  wire [3:0]DDR_dqs_n;
  wire [3:0]DDR_dqs_p;
  wire DDR_odt;
  wire DDR_ras_n;
  wire DDR_reset_n;
  wire DDR_we_n;
  wire FIXED_IO_ddr_vrn;
  wire FIXED_IO_ddr_vrp;
  wire [53:0]FIXED_IO_mio;
  wire FIXED_IO_ps_clk;
  wire FIXED_IO_ps_porb;
  wire FIXED_IO_ps_srstb;
  wire GMII_ETHERNET_1_col;
  wire GMII_ETHERNET_1_crs;
  wire GMII_ETHERNET_1_rx_clk;
  wire GMII_ETHERNET_1_rx_dv;
  wire GMII_ETHERNET_1_rx_er;
  wire [7:0]GMII_ETHERNET_1_rxd;
  wire GMII_ETHERNET_1_tx_clk;
  wire [0:0]GMII_ETHERNET_1_tx_en;
  wire [0:0]GMII_ETHERNET_1_tx_er;
  wire [7:0]GMII_ETHERNET_1_txd;
  wire [0:0]btns_5bits_tri_i_0;
  wire [1:1]btns_5bits_tri_i_1;
  wire [2:2]btns_5bits_tri_i_2;
  wire [3:3]btns_5bits_tri_i_3;
  wire [4:4]btns_5bits_tri_i_4;
  wire [0:0]btns_5bits_tri_io_0;
  wire [1:1]btns_5bits_tri_io_1;
  wire [2:2]btns_5bits_tri_io_2;
  wire [3:3]btns_5bits_tri_io_3;
  wire [4:4]btns_5bits_tri_io_4;
  wire [0:0]btns_5bits_tri_o_0;
  wire [1:1]btns_5bits_tri_o_1;
  wire [2:2]btns_5bits_tri_o_2;
  wire [3:3]btns_5bits_tri_o_3;
  wire [4:4]btns_5bits_tri_o_4;
  wire [0:0]btns_5bits_tri_t_0;
  wire [1:1]btns_5bits_tri_t_1;
  wire [2:2]btns_5bits_tri_t_2;
  wire [3:3]btns_5bits_tri_t_3;
  wire [4:4]btns_5bits_tri_t_4;
  wire [7:0]leds_8bits_tri_o;

IOBUF btns_5bits_tri_iobuf_0
       (.I(btns_5bits_tri_o_0),
        .IO(btns_5bits_tri_io[0]),
        .O(btns_5bits_tri_i_0),
        .T(btns_5bits_tri_t_0));
IOBUF btns_5bits_tri_iobuf_1
       (.I(btns_5bits_tri_o_1),
        .IO(btns_5bits_tri_io[1]),
        .O(btns_5bits_tri_i_1),
        .T(btns_5bits_tri_t_1));
IOBUF btns_5bits_tri_iobuf_2
       (.I(btns_5bits_tri_o_2),
        .IO(btns_5bits_tri_io[2]),
        .O(btns_5bits_tri_i_2),
        .T(btns_5bits_tri_t_2));
IOBUF btns_5bits_tri_iobuf_3
       (.I(btns_5bits_tri_o_3),
        .IO(btns_5bits_tri_io[3]),
        .O(btns_5bits_tri_i_3),
        .T(btns_5bits_tri_t_3));
IOBUF btns_5bits_tri_iobuf_4
       (.I(btns_5bits_tri_o_4),
        .IO(btns_5bits_tri_io[4]),
        .O(btns_5bits_tri_i_4),
        .T(btns_5bits_tri_t_4));
pfSenseZ pfSenseZ_i
       (.DDR_addr(DDR_addr),
        .DDR_ba(DDR_ba),
        .DDR_cas_n(DDR_cas_n),
        .DDR_ck_n(DDR_ck_n),
        .DDR_ck_p(DDR_ck_p),
        .DDR_cke(DDR_cke),
        .DDR_cs_n(DDR_cs_n),
        .DDR_dm(DDR_dm),
        .DDR_dq(DDR_dq),
        .DDR_dqs_n(DDR_dqs_n),
        .DDR_dqs_p(DDR_dqs_p),
        .DDR_odt(DDR_odt),
        .DDR_ras_n(DDR_ras_n),
        .DDR_reset_n(DDR_reset_n),
        .DDR_we_n(DDR_we_n),
        .FIXED_IO_ddr_vrn(FIXED_IO_ddr_vrn),
        .FIXED_IO_ddr_vrp(FIXED_IO_ddr_vrp),
        .FIXED_IO_mio(FIXED_IO_mio),
        .FIXED_IO_ps_clk(FIXED_IO_ps_clk),
        .FIXED_IO_ps_porb(FIXED_IO_ps_porb),
        .FIXED_IO_ps_srstb(FIXED_IO_ps_srstb),
        .GMII_ETHERNET_1_col(GMII_ETHERNET_1_col),
        .GMII_ETHERNET_1_crs(GMII_ETHERNET_1_crs),
        .GMII_ETHERNET_1_rx_clk(GMII_ETHERNET_1_rx_clk),
        .GMII_ETHERNET_1_rx_dv(GMII_ETHERNET_1_rx_dv),
        .GMII_ETHERNET_1_rx_er(GMII_ETHERNET_1_rx_er),
        .GMII_ETHERNET_1_rxd(GMII_ETHERNET_1_rxd),
        .GMII_ETHERNET_1_tx_clk(GMII_ETHERNET_1_tx_clk),
        .GMII_ETHERNET_1_tx_en(GMII_ETHERNET_1_tx_en),
        .GMII_ETHERNET_1_tx_er(GMII_ETHERNET_1_tx_er),
        .GMII_ETHERNET_1_txd(GMII_ETHERNET_1_txd),
        .btns_5bits_tri_i({btns_5bits_tri_i_4,btns_5bits_tri_i_3,btns_5bits_tri_i_2,btns_5bits_tri_i_1,btns_5bits_tri_i_0}),
        .btns_5bits_tri_o({btns_5bits_tri_o_4,btns_5bits_tri_o_3,btns_5bits_tri_o_2,btns_5bits_tri_o_1,btns_5bits_tri_o_0}),
        .btns_5bits_tri_t({btns_5bits_tri_t_4,btns_5bits_tri_t_3,btns_5bits_tri_t_2,btns_5bits_tri_t_1,btns_5bits_tri_t_0}),
        .leds_8bits_tri_o(leds_8bits_tri_o));
endmodule
